--------------------------------------------------------------------------------
-- Project    : <project title> 
--------------------------------------------------------------------------------
-- File       : <filename> 
-- Author     : Kelve T. Henrique
-- Company    : FH Technikum Wien
-- Last update: <date> 
-- Platform   : Linux, ModelSim, Xilinx Vivado
--------------------------------------------------------------------------------
-- Description: <What is this code for?> 
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all; -- use logic elements
