---------------------------------------------------------------------------- 
--  <PROJECT TITLE> - <BEGINNING DATE>
----------------------------------------------------------------------------
--! @file <file_name>
--! @author Kelve T. Henrique
--! @date dd Mmm, YYYY
--! @version 1.0
--!
--! @brief   <What is this code>
--!
--! @details <Description of what is gonna be done here>
----------------------------------------------------------------------------

